`timescale 10ps/10ps

module instructionFetch (clk, reset, instruction, currentPC, branchAddress, brTaken);