/*	3:8 Decoder. Building block of 5:32 decoder - regDecoder
 * Depending on the en signal, it will choose what to output
 *	Input: en, [2:0] in
 * Output: [7:0] out
 */
`timescale 1ns/10ps
